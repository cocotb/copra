package multi_dim_array_pkg;

    typedef logic               [2:0] test_array_entry_t;
    typedef test_array_entry_t  [2:0] test_2d_array_t;
    typedef test_2d_array_t     [2:0] test_3d_array_t;

endpackage 
